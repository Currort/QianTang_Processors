module ID(
    input               clk_sys_i      ,
    input [31:0] instr_i,
    output [31:0] rst1,
    output [31:0] rst2,
    output [31:0] rd,

);
    always @(posedge clk_sys_i) begin
        ;
    end

endmodule //ID
