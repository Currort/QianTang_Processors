module PC
#(
    localparam ADDR_WIDTH =  'd16
)(
    input   clk_sys_i   ,     
    input  [31:0] iaddr_i     ,     
    input  add4_en_i , 
    input  
    output [31:0] iaddr_o
);
    

endmodule //PC

